LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY hw_image_generator IS
  GENERIC(
    pixels_y :  INTEGER := 478;   -- row that first color will persist until
    pixels_x :  INTEGER := 600     -- column that first color will persist until
  );
  PORT(
    disp_ena :  IN   STD_LOGIC;  -- display enable ('1' = display time, '0' = blanking time)
    row      :  IN   INTEGER;    -- row pixel coordinate
    column   :  IN   INTEGER;    -- column pixel coordinate
    red      :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');  -- red magnitude output to DAC
    green    :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');  -- green magnitude output to DAC
    blue     :  OUT  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0')   -- blue magnitude output to DAC
  );
END hw_image_generator;

ARCHITECTURE behavior OF hw_image_generator IS

  -- Character 'S' bitmap in 20x100 format, each bit represents a 20x20 block
  TYPE bitmap_array IS ARRAY (0 TO 19) OF STD_LOGIC_VECTOR(99 DOWNTO 0);
  CONSTANT char_S : bitmap_array := (
    "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", 
    "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
    "0001000000001000111111111000001111111110011111111100100000000010000000000101111111100111111110000000",
    "0001000000001000000010000000001000000010010000000100100000000010000000000100000000100100000000000000",
    "0001000000001000000010000000001000000010010000000100100000000010000000000100000000100100000000000000",
    "0001000000001000000010000000001000000010010000000100100000000010000000000100000000100100000000000000",
    "0001000000001000000010000000001000000010011111111100100000000010000000000101111111100100000000000000",
    "0001000000001000000010000000001000000010010000000100100000000010000000000100000000100111111110000000",
    "0001000000001000000010000000001000000010010000000100100000000010000000000100000000100000000010000000",
    "0001000000001000000010000000001000000010010000000100100000000010000000000100000000100000000010000000",
    "0001000000001000000010000000001000000010010000000100100000000010000000000100000000100000000010000000", 
    "0001111111111000000010000000001111111110010000000100111111110011111111100100000000100111111110000000", 
    "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", 
    "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", 
    "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", 
    "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", 
    "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", 
    "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", 
    "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000", 
    "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"  
  );

BEGIN
  PROCESS(disp_ena, row, column)
  BEGIN

    IF (disp_ena = '1') THEN  -- display time
      -- Set the background to white
      red <= (OTHERS => '1');    
      green <= (OTHERS => '1');  
      blue <= (OTHERS => '1');   

-- Assuming char_S is a 20x100 array of std_logic representing the character bitmap
-- This example assumes char_S is declared as follows:
-- type char_array is array (0 to 19) of std_logic_vector(99 downto 0);
-- signal char_S : char_array;

-- Loop through the character bitmap for "S"
    FOR i IN 0 TO 19 LOOP  -- 20 rows (flipped)
    IF (row >= (450 + i * 10) AND row < (470 + i * 10)) THEN  -- Scale rows by 10
        FOR j IN 0 TO 99 LOOP  -- 100 columns
            IF (column >= (550 + j * 10) AND column < (570 + j * 10)) THEN  -- Scale columns by 10
                IF (char_S(i)(99 - j) = '1') THEN  -- Flip the bitmap horizontally
                    -- Set pixel color to black for "S"
                    red <= X"FF";   -- Assign all bits to '0'
                    green <= X"A5"; -- Assign all bits to '0'
                    blue <=  X"00";  -- Assign all bits to '0'
                END IF;
            END IF;
        END LOOP;
    END IF;
END LOOP;




    ELSE  -- blanking time
      red <= (OTHERS => '0');
      green <= (OTHERS => '0');
      blue <= (OTHERS => '0');
    END IF;

  END PROCESS;
END behavior;
